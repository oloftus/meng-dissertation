library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

package Constants is
    constant precisionConst : INTEGER := 8;
end package Constants;
